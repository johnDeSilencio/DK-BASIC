module gamecube_bit_decoder (
    input CLK,
    input n_RST,
    input DIR,
    input n_SEND,
    input TO_GAMECUBE,
    output reg DATALINE,
    output reg FROM_GAMECUBE,
    output reg BUSY,
    output reg LOAD
);
    reg 
endmodule